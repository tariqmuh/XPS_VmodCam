library verilog;
use verilog.vl_types.all;
entity user_logic is
    generic(
        HDMI_HRES       : integer := 640;
        HDMI_BYTES_PER_PIXEL: integer := 4;
        C_MST_NATIVE_DATA_WIDTH: integer := 32;
        C_LENGTH_WIDTH  : integer := 12;
        C_MST_AWIDTH    : integer := 32;
        C_NUM_REG       : integer := 4;
        C_SLV_DWIDTH    : integer := 32;
        CMD_IDLE        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        CMD_RUN         : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        CMD_WAIT_FOR_DATA: vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        CMD_DONE        : vl_logic_vector(1 downto 0) := (Hi1, Hi1);
        LLRD_IDLE       : vl_logic := Hi0;
        LLRD_GO         : vl_logic := Hi1;
        LLWR_IDLE       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        LLWR_SNGL_INIT  : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        LLWR_SNGL       : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        LLWR_BRST_INIT  : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        LLWR_BRST       : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        LLWR_BRST_LAST_BEAT: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        BE_WIDTH        : vl_notype;
        BYTES_PER_BEAT  : vl_notype;
        GO_DATA_KEY     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        GO_BYTE_LANE    : integer := 15
    );
    port(
        PXL_CLK_X1      : in     vl_logic;
        PXL_CLK_X2      : in     vl_logic;
        PXL_CLK_X10     : in     vl_logic;
        PXL_PLL_LOCKED  : in     vl_logic;
        TMDS            : out    vl_logic_vector(3 downto 0);
        TMDSB           : out    vl_logic_vector(3 downto 0);
        Bus2IP_Clk      : in     vl_logic;
        Bus2IP_Resetn   : in     vl_logic;
        Bus2IP_Data     : in     vl_logic_vector;
        Bus2IP_BE       : in     vl_logic_vector;
        Bus2IP_RdCE     : in     vl_logic_vector;
        Bus2IP_WrCE     : in     vl_logic_vector;
        IP2Bus_Data     : out    vl_logic_vector;
        IP2Bus_RdAck    : out    vl_logic;
        IP2Bus_WrAck    : out    vl_logic;
        IP2Bus_Error    : out    vl_logic;
        ip2bus_mstrd_req: out    vl_logic;
        ip2bus_mstwr_req: out    vl_logic;
        ip2bus_mst_addr : out    vl_logic_vector;
        ip2bus_mst_be   : out    vl_logic_vector;
        ip2bus_mst_length: out    vl_logic_vector;
        ip2bus_mst_type : out    vl_logic;
        ip2bus_mst_lock : out    vl_logic;
        ip2bus_mst_reset: out    vl_logic;
        bus2ip_mst_cmdack: in     vl_logic;
        bus2ip_mst_cmplt: in     vl_logic;
        bus2ip_mst_error: in     vl_logic;
        bus2ip_mst_rearbitrate: in     vl_logic;
        bus2ip_mst_cmd_timeout: in     vl_logic;
        bus2ip_mstrd_d  : in     vl_logic_vector;
        bus2ip_mstrd_rem: in     vl_logic_vector;
        bus2ip_mstrd_sof_n: in     vl_logic;
        bus2ip_mstrd_eof_n: in     vl_logic;
        bus2ip_mstrd_src_rdy_n: in     vl_logic;
        bus2ip_mstrd_src_dsc_n: in     vl_logic;
        ip2bus_mstrd_dst_rdy_n: out    vl_logic;
        ip2bus_mstrd_dst_dsc_n: out    vl_logic;
        ip2bus_mstwr_d  : out    vl_logic_vector;
        ip2bus_mstwr_rem: out    vl_logic_vector;
        ip2bus_mstwr_src_rdy_n: out    vl_logic;
        ip2bus_mstwr_src_dsc_n: out    vl_logic;
        ip2bus_mstwr_sof_n: out    vl_logic;
        ip2bus_mstwr_eof_n: out    vl_logic;
        bus2ip_mstwr_dst_rdy_n: in     vl_logic;
        bus2ip_mstwr_dst_dsc_n: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of HDMI_HRES : constant is 1;
    attribute mti_svvh_generic_type of HDMI_BYTES_PER_PIXEL : constant is 1;
    attribute mti_svvh_generic_type of C_MST_NATIVE_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_LENGTH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_MST_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_NUM_REG : constant is 1;
    attribute mti_svvh_generic_type of C_SLV_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of CMD_IDLE : constant is 2;
    attribute mti_svvh_generic_type of CMD_RUN : constant is 2;
    attribute mti_svvh_generic_type of CMD_WAIT_FOR_DATA : constant is 2;
    attribute mti_svvh_generic_type of CMD_DONE : constant is 2;
    attribute mti_svvh_generic_type of LLRD_IDLE : constant is 1;
    attribute mti_svvh_generic_type of LLRD_GO : constant is 1;
    attribute mti_svvh_generic_type of LLWR_IDLE : constant is 2;
    attribute mti_svvh_generic_type of LLWR_SNGL_INIT : constant is 2;
    attribute mti_svvh_generic_type of LLWR_SNGL : constant is 2;
    attribute mti_svvh_generic_type of LLWR_BRST_INIT : constant is 2;
    attribute mti_svvh_generic_type of LLWR_BRST : constant is 2;
    attribute mti_svvh_generic_type of LLWR_BRST_LAST_BEAT : constant is 2;
    attribute mti_svvh_generic_type of BE_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of BYTES_PER_BEAT : constant is 3;
    attribute mti_svvh_generic_type of GO_DATA_KEY : constant is 2;
    attribute mti_svvh_generic_type of GO_BYTE_LANE : constant is 1;
end user_logic;
